entity hello_world is
end entity;

architecture sim of hello_world is
begin
	process is
	begin
		report "hello world!!!!!333433444";
		wait;
	
	end process;
end architecture;